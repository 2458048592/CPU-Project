`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:10:47 08/26/2015 
// Design Name: 
// Module Name:    font_table 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module font_table(
			input wire [7:0] ascii,
			input wire [9:0] font_address,
			output font_dot
    );

	parameter font = {
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h0000000000000000,
			64'h1818181800181800,
			64'h6c6c480000000000,
			64'h6c6cfe6cfe6c6c00,
			64'h187ed87e1b7e1800,
			64'h62660c1830664600,
			64'h386c6876dccc7600,
			64'h1818300000000000,
			64'h0c18303030180c00,
			64'h30180c0c0c183000,
			64'h006c38fe386c0000,
			64'h0018187e18180000,
			64'h0000000000181810,
			64'h0000007e00000000,
			64'h0000000000181800,
			64'h02060c1830604000,
			64'h3c666e7666663c00,
			64'h1818381818183c00,
			64'h7c06063c60607c00,
			64'h7c06063c06067c00,
			64'h6666667e06060600,
			64'h7e60607c06067c00,
			64'h3c60607c66663c00,
			64'h7e060c1818181800,
			64'h3c66663c66663c00,
			64'h3c66663e06063c00,
			64'h0018180018180000,
			64'h0000181800181810,
			64'h0c18306030180c00,
			64'h00007e007e000000,
			64'h30180c060c183000,
			64'h3c66061c18001800,
			64'h3c666e6a6e603e00,
			64'h3c66667e66666600,
			64'h7c66667c66667c00,
			64'h3c66606060663c00,
			64'h7c66666666667c00,
			64'h7e60607c60607e00,
			64'h7e60607c60606000,
			64'h3c66606e66663c00,
			64'h6666667e66666600,
			64'h3c18181818183c00,
			64'h3e0c0c0c0c6c3800,
			64'h666c7870786c6600,
			64'h6060606060607e00,
			64'hc6eefed6c6c6c600,
			64'h6666767e6e666600,
			64'h3c66666666663c00,
			64'h7c66667c60606000,
			64'h3c6666666e663e00,
			64'h7c66667c66666600,
			64'h3e60603c06067c00,
			64'h7e18181818181800,
			64'h6666666666663c00,
			64'h666666663c3c1800,
			64'hc6c6d6d6feee4400,
			64'h66663c183c666600,
			64'h6666663c18181800,
			64'h7e060c1830607e00,
			64'h3c30303030303c00,
			64'h406030180c060200,
			64'h3c0c0c0c0c0c3c00,
			64'h10386c0000000000,
			64'h00000000000000ff,
			64'h18180c0000000000,
			64'h00003c063e663a00,
			64'h60607c6666667c00,
			64'h00003c6660663c00,
			64'h06063e6666663e00,
			64'h00003c667c603c00,
			64'h0e18183e18181800,
			64'h00003e66663e063c,
			64'h60607c6666666600,
			64'h1800181818181800,
			64'h1800181818181870,
			64'h6060666c786c6600,
			64'h3030303030301c00,
			64'h0000ccfed6c6c600,
			64'h00007c6666666600,
			64'h00003c6666663c00,
			64'h00007c66667c6060,
			64'h00003e66663e0606,
			64'h0000363830303000,
			64'h00003e603c067c00,
			64'h18183c1818180c00,
			64'h0000666666663c00,
			64'h00006666663c1800,
			64'h0000c6d6d67c2800,
			64'h0000663c183c6600,
			64'h00006666663e067c,
			64'h00007e0c18307e00,
			64'h1c30306030301c00,
			64'h1818181818181800,
			64'h380c0c060c0c3800,
			64'h00324c0000000000,
			64'h0000000000000000
	};

	assign font_dot = font[(127 - ascii)*64 + 63 - font_address];

endmodule
